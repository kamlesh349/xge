`include "uvm.sv"
`include "uvm_macros.svh"
import uvm_pkg::*;

`include "rx_env.sv"
`include "my_test.sv"
`include "top.sv"
