`include   "uvm_macros.svh"
 import     uvm_pkg::*;

`include   "xge_ifc.sv"
`include"agent/header.svh"
`include "env.sv"
`include "test.sv"
`include "top.sv"
