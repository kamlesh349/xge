class xge_mon extends uvm_monitor;
	`uvm_componet_utils(xge_mon)
	vxge		vif;
	xge_pkt	rx,tx;

	uvm_analysis_port#(xge_pkt)	nq_ap;

	function new(string name="xge_mon", uvm_componet parent);
		super.new(name, parent);
		nq_ap = new("nq_ap",this);
	endfunction

	function void build_phase(uvm_phase phase);
		if (!uvm_config_db#(vif)::get(this,"","xge_ifc",vif)
			`uvm_fatal("MON", "failed to get interface")
	endfunction

	task run_phase(uvm_phase phase);
		forever begin
			tx	= xge_pkt::type_id::create("tx",this);
			rx	= xge_pkt::type_id::create("rx",this);
		fork
			begin:  rst
				wait(!vif.reset_156m25_n);
				`uvm_info(get_type_name(),"_Reset_applied",UVM_MEDIUM)
				dq_ap.write(rx);
				nq_ap.write(tx);
				disable rx_dq
				disable tx_nq
				while(!vif.reset_156m25_n);
			end:    rst
			begin:  tx_dq
				wait(vif.cbtxrx.pkt_tx_sop);
				do begin
					tx.data.push_back(vif.cbtxrx.pkt_tx_data);
					@(vif.cbtxrx);
				end while(!vif.cbtxrx.pkt_tx_eop);
				tx.data.push_back(vif.cbtxrx.pkt_tx_data);
				$cast(tx.mod, vif.cbtxrx.pkt_tx_mod);
			end:    tx_dq
			begin:  rx_nq
				wait(vif.cbtxrx.pkt_rx_sop);
				do begin
					rx.data.push_back(vif.cbtxrx.pkt_rx_data);
					@(vif.cbtxrx);
				end while(!vif.cbtxrx.pkt_rx_eop);
				rx.data.push_back(vif.cbtxrx.pkt_rx_data);
				$cast(rx.mod, vif.cbtxrx.pkt_rx_mod);
			end:    rx_nq
		join_any
		end//4ever
	endtask
endclass
